module fetchstage0_tb;
endmodule