module memorystage1_tb;
endmodule
