`ifndef BUSINTERFACE_H

localparam  CW_LONG = 2'b00,
            CW_WORD = 2'b01,
            CW_BYTE = 2'b10,
            CW_NULL = 2'b11;

`define BUSINTERFACE_H 1
`endif
