`ifndef REGISTERS_VH

// Imediate write types
localparam  IT_TOP = 2'b00,
            IT_BOTTOM = 2'b01,
            IT_UNSIGNED = 2'b10,
            IT_SIGNED = 2'b11;

`define REGISTERS_VH 1
`endif
