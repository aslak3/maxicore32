typedef reg [4:0] t_opcode;

localparam t_opcode OPCODE_NOP      = 5'b00000;
