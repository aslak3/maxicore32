`ifndef REGISTERS_VH
typedef reg [31:0] t_reg;
typedef t_reg t_regs [16];
typedef reg [3:0] t_reg_index;

`define REGISTERS_VH 1
`endif
