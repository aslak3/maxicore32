module registersstage2_tb;
endmodule
