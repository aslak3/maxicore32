typedef reg [4:0] t_alu_op;
